`timescale 1ns/1ns
`include "q1ha.v"

module q1ha_tb();
reg x,y;
wire sum, c_out;

q1ha l4(x,y,sum, c_out);
initial
begin

  $dumpfile("q1ha_tb.vcd");
  $dumpvars(0, q1ha_tb);
  
  x=1'b0; y=1'b0; 
  #20;
  
  x=1'b0; y=1'b1;
  #20;
  
  x=1'b1; y=1'b0; 
  #20;

  x=1'b1; y=1'b1; 
  #20;

   $display("test complete");
end 

endmodule
